module encoder (
  input [15:0] in,
  output reg [3:0] out
);

always @(*) begin
  case (in)
    16'b0000_0000_0000_0001: out = 4'b0000; // 0
    16'b0000_0000_0000_0010: out = 4'b0001; // 1
    16'b0000_0000_0000_0100: out = 4'b0010; // 2
    16'b0000_0000_0000_1000: out = 4'b0011; // 3
    16'b0000_0000_0001_0000: out = 4'b0100; // 4
    16'b0000_0000_0010_0000: out = 4'b0101; // 5
    16'b0000_0000_0100_0000: out = 4'b0110; // 6
    16'b0000_0000_1000_0000: out = 4'b0111; // 7
    16'b0000_0001_0000_0000: out = 4'b1000; // 8
    16'b0000_0010_0000_0000: out = 4'b1001; // 9
    16'b0000_0100_0000_0000: out = 4'b1010; // 10
    16'b0000_1000_0000_0000: out = 4'b1011; // 11
    16'b0001_0000_0000_0000: out = 4'b1100; // 12
    16'b0010_0000_0000_0000: out = 4'b1101; // 13
    16'b0100_0000_0000_0000: out = 4'b1110; // 14
    16'b1000_0000_0000_0000: out = 4'b1111; // 15
    default: out = 4'bxxxx; 
  endcase
end

endmodule
